module alu_less_than(
    input logic [31:0]      i_a,
    input logic [31:0]      i_b,
    input logic             sign,   // 1: unsign, 0 sign
    output logic [31:0]     o_slt
);



endmodule
